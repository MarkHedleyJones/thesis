electrodeModel
****************************************
*        Faradaic branch start         *
****************************************
.SUBCKT faradaic n1 n2
.PARAM Vt=0.025875
.PARAM i0=2.75674884748e-12
.PARAM n=1.35992195766
.PARAM nVt=n*Vt
Bdm1 n1 n2 I=i0*exp(v(n1,n2)/nVt)
Bdm2 n2 n1 I=i0*exp(v(n2,n1)/nVt)
R_b n1 n2 1e10
.ENDS faradaic
****************************************
*         Resistor ladder start        *
****************************************
.SUBCKT ladder e1 e2 e3 e4 e5 e6 e7 e8
RRAD_1_1 1 2 24.2043775561
RRAD_1_2 2 3 24.2043775561
RRAD_1_3 3 4 24.2043775561
RRAD_1_4 4 5 24.2043775561
RRAD_1_5 5 1000 24.2043775561
RVERT_2_1 1 6 220.634498116
RVERT_2_2 2 7 55.158624529
RVERT_2_3 3 8 13.7896561322
RVERT_2_4 4 9 3.44741403306
RVERT_2_5 5 10 0.861853508265
RRAD_3_1 6 7 24.2043775561
RRAD_3_2 7 8 24.2043775561
RRAD_3_3 8 9 24.2043775561
RRAD_3_4 9 10 24.2043775561
RRAD_3_5 10 1000 24.2043775561
RVERT_4_1 6 11 220.634498116
RVERT_4_2 7 12 55.158624529
RVERT_4_3 8 13 13.7896561322
RVERT_4_4 9 14 3.44741403306
RVERT_4_5 10 15 0.861853508265
RRAD_5_1 11 12 24.2043775561
RRAD_5_2 12 13 24.2043775561
RRAD_5_3 13 14 24.2043775561
RRAD_5_4 14 15 24.2043775561
RRAD_5_5 15 1000 24.2043775561
RVERT_6_1 11 e1 220.634498116
RVERT_6_2 12 17 55.158624529
RVERT_6_3 13 18 13.7896561322
RVERT_6_4 14 19 3.44741403306
RVERT_6_5 15 20 0.861853508265
RRAD_7_1 e1 17 24.2043775561
RRAD_7_2 17 18 24.2043775561
RRAD_7_3 18 19 24.2043775561
RRAD_7_4 19 20 24.2043775561
RRAD_7_5 20 1000 24.2043775561
RVERT_8_1 e1 21 220.634498116
RVERT_8_2 17 22 55.158624529
RVERT_8_3 18 23 13.7896561322
RVERT_8_4 19 24 3.44741403306
RVERT_8_5 20 25 0.861853508265
RRAD_9_1 21 22 18.1532831671
RRAD_9_2 22 23 18.1532831671
RRAD_9_3 23 24 18.1532831671
RRAD_9_4 24 25 18.1532831671
RRAD_9_5 25 1000 18.1532831671
RVERT_10_1 21 e2 220.634498116
RVERT_10_2 22 27 55.158624529
RVERT_10_3 23 28 13.7896561322
RVERT_10_4 24 29 3.44741403306
RVERT_10_5 25 30 0.861853508265
RRAD_11_1 e2 27 24.2043775561
RRAD_11_2 27 28 24.2043775561
RRAD_11_3 28 29 24.2043775561
RRAD_11_4 29 30 24.2043775561
RRAD_11_5 30 1000 24.2043775561
RVERT_12_1 e2 31 220.634498116
RVERT_12_2 27 32 55.158624529
RVERT_12_3 28 33 13.7896561322
RVERT_12_4 29 34 3.44741403306
RVERT_12_5 30 35 0.861853508265
RRAD_13_1 31 32 18.1532831671
RRAD_13_2 32 33 18.1532831671
RRAD_13_3 33 34 18.1532831671
RRAD_13_4 34 35 18.1532831671
RRAD_13_5 35 1000 18.1532831671
RVERT_14_1 31 e3 220.634498116
RVERT_14_2 32 37 55.158624529
RVERT_14_3 33 38 13.7896561322
RVERT_14_4 34 39 3.44741403306
RVERT_14_5 35 40 0.861853508265
RRAD_15_1 e3 37 24.2043775561
RRAD_15_2 37 38 24.2043775561
RRAD_15_3 38 39 24.2043775561
RRAD_15_4 39 40 24.2043775561
RRAD_15_5 40 1000 24.2043775561
RVERT_16_1 e3 41 220.634498116
RVERT_16_2 37 42 55.158624529
RVERT_16_3 38 43 13.7896561322
RVERT_16_4 39 44 3.44741403306
RVERT_16_5 40 45 0.861853508265
RRAD_17_1 41 42 18.1532831671
RRAD_17_2 42 43 18.1532831671
RRAD_17_3 43 44 18.1532831671
RRAD_17_4 44 45 18.1532831671
RRAD_17_5 45 1000 18.1532831671
RVERT_18_1 41 e4 220.634498116
RVERT_18_2 42 47 55.158624529
RVERT_18_3 43 48 13.7896561322
RVERT_18_4 44 49 3.44741403306
RVERT_18_5 45 50 0.861853508265
RRAD_19_1 e4 47 24.2043775561
RRAD_19_2 47 48 24.2043775561
RRAD_19_3 48 49 24.2043775561
RRAD_19_4 49 50 24.2043775561
RRAD_19_5 50 1000 24.2043775561
RVERT_20_1 e4 51 220.634498116
RVERT_20_2 47 52 55.158624529
RVERT_20_3 48 53 13.7896561322
RVERT_20_4 49 54 3.44741403306
RVERT_20_5 50 55 0.861853508265
RRAD_21_1 51 52 18.1532831671
RRAD_21_2 52 53 18.1532831671
RRAD_21_3 53 54 18.1532831671
RRAD_21_4 54 55 18.1532831671
RRAD_21_5 55 1000 18.1532831671
RVERT_22_1 51 e5 220.634498116
RVERT_22_2 52 57 55.158624529
RVERT_22_3 53 58 13.7896561322
RVERT_22_4 54 59 3.44741403306
RVERT_22_5 55 60 0.861853508265
RRAD_23_1 e5 57 24.2043775561
RRAD_23_2 57 58 24.2043775561
RRAD_23_3 58 59 24.2043775561
RRAD_23_4 59 60 24.2043775561
RRAD_23_5 60 1000 24.2043775561
RVERT_24_1 e5 61 220.634498116
RVERT_24_2 57 62 55.158624529
RVERT_24_3 58 63 13.7896561322
RVERT_24_4 59 64 3.44741403306
RVERT_24_5 60 65 0.861853508265
RRAD_25_1 61 62 18.1532831671
RRAD_25_2 62 63 18.1532831671
RRAD_25_3 63 64 18.1532831671
RRAD_25_4 64 65 18.1532831671
RRAD_25_5 65 1000 18.1532831671
RVERT_26_1 61 e6 220.634498116
RVERT_26_2 62 67 55.158624529
RVERT_26_3 63 68 13.7896561322
RVERT_26_4 64 69 3.44741403306
RVERT_26_5 65 70 0.861853508265
RRAD_27_1 e6 67 24.2043775561
RRAD_27_2 67 68 24.2043775561
RRAD_27_3 68 69 24.2043775561
RRAD_27_4 69 70 24.2043775561
RRAD_27_5 70 1000 24.2043775561
RVERT_28_1 e6 71 220.634498116
RVERT_28_2 67 72 55.158624529
RVERT_28_3 68 73 13.7896561322
RVERT_28_4 69 74 3.44741403306
RVERT_28_5 70 75 0.861853508265
RRAD_29_1 71 72 18.1532831671
RRAD_29_2 72 73 18.1532831671
RRAD_29_3 73 74 18.1532831671
RRAD_29_4 74 75 18.1532831671
RRAD_29_5 75 1000 18.1532831671
RVERT_30_1 71 e7 220.634498116
RVERT_30_2 72 77 55.158624529
RVERT_30_3 73 78 13.7896561322
RVERT_30_4 74 79 3.44741403306
RVERT_30_5 75 80 0.861853508265
RRAD_31_1 e7 77 24.2043775561
RRAD_31_2 77 78 24.2043775561
RRAD_31_3 78 79 24.2043775561
RRAD_31_4 79 80 24.2043775561
RRAD_31_5 80 1000 24.2043775561
RVERT_32_1 e7 81 220.634498116
RVERT_32_2 77 82 55.158624529
RVERT_32_3 78 83 13.7896561322
RVERT_32_4 79 84 3.44741403306
RVERT_32_5 80 85 0.861853508265
RRAD_33_1 81 82 18.1532831671
RRAD_33_2 82 83 18.1532831671
RRAD_33_3 83 84 18.1532831671
RRAD_33_4 84 85 18.1532831671
RRAD_33_5 85 1000 18.1532831671
RVERT_34_1 81 e8 220.634498116
RVERT_34_2 82 87 55.158624529
RVERT_34_3 83 88 13.7896561322
RVERT_34_4 84 89 3.44741403306
RVERT_34_5 85 90 0.861853508265
RRAD_35_1 e8 87 24.2043775561
RRAD_35_2 87 88 24.2043775561
RRAD_35_3 88 89 24.2043775561
RRAD_35_4 89 90 24.2043775561
RRAD_35_5 90 1000 24.2043775561
RVERT_36_1 e8 91 220.634498116
RVERT_36_2 87 92 55.158624529
RVERT_36_3 88 93 13.7896561322
RVERT_36_4 89 94 3.44741403306
RVERT_36_5 90 95 0.861853508265
RRAD_37_1 91 92 24.2043775561
RRAD_37_2 92 93 24.2043775561
RRAD_37_3 93 94 24.2043775561
RRAD_37_4 94 95 24.2043775561
RRAD_37_5 95 1000 24.2043775561
RVERT_38_1 91 96 220.634498116
RVERT_38_2 92 97 55.158624529
RVERT_38_3 93 98 13.7896561322
RVERT_38_4 94 99 3.44741403306
RVERT_38_5 95 100 0.861853508265
RRAD_39_1 96 97 24.2043775561
RRAD_39_2 97 98 24.2043775561
RRAD_39_3 98 99 24.2043775561
RRAD_39_4 99 100 24.2043775561
RRAD_39_5 100 1000 24.2043775561
RVERT_40_1 96 101 220.634498116
RVERT_40_2 97 102 55.158624529
RVERT_40_3 98 103 13.7896561322
RVERT_40_4 99 104 3.44741403306
RVERT_40_5 100 105 0.861853508265
RRAD_41_1 101 102 24.2043775561
RRAD_41_2 102 103 24.2043775561
RRAD_41_3 103 104 24.2043775561
RRAD_41_4 104 105 24.2043775561
RRAD_41_5 105 1000 24.2043775561
.ENDS ladder
****************************************
*           Fracpole/CPE start         *
****************************************
.SUBCKT displacement a b
R0 a 1 42769491660.0
C0 1 b 0.000359405061629
R1 a 2 23314469349.4
C1 2 b 0.00030602676341
R2 a 3 12709163937.9
C2 3 b 0.000260576129615
R3 a 4 6928008764.81
C3 4 b 0.000221875755469
R4 a 5 3776590315.45
C4 5 b 0.000188923102579
R5 a 6 2058691738.85
C5 6 b 0.000160864528044
R6 a 7 1122232310.52
C6 7 b 0.000136973170722
R7 a 8 611750333.967
C7 8 b 0.000116630121791
R8 a 9 333476827.926
C8 9 b 9.93083918356e-05
R9 a 10 181784608.179
C9 10 b 8.45592591134e-05
R10 a 11 99094272.8358
C10 11 b 7.20006453598e-05
R11 a 12 54018186.7277
C11 12 b 6.13072179982e-05
R12 a 13 29446348.5512
C12 13 b 5.22019623559e-05
R13 a 14 16051768.775
C13 14 b 4.44490055623e-05
R14 a 15 8750126.70443
C14 15 b 3.78475062299e-05
R15 a 16 4769861.71536
C15 16 b 3.22264516315e-05
R16 a 17 2600143.0096
C16 17 b 2.74402275925e-05
R17 a 18 1417387.77219
C17 18 b 2.33648463361e-05
R18 a 19 772645.231177
C18 19 b 1.98947345633e-05
R19 a 20 421183.719075
C19 20 b 1.69399985624e-05
R20 a 21 229595.314972
C20 21 b 1.44240955003e-05
R21 a 22 125156.805142
C21 22 b 1.22818505702e-05
R22 a 23 68225.3724348
C22 23 b 1.04577686292e-05
R23 a 24 37190.9576838
C23 24 b 8.90459658967e-06
R24 a 25 20273.5035967
C24 25 b 7.5820993212e-06
R25 a 26 11051.4752424
C25 26 b 6.45601735437e-06
R26 a 27 6024.37089629
C26 27 b 5.49717938452e-06
R27 a 28 3284.0
C27 28 b 4.68074658522e-06
R28 a 29 1790.17132007
C28 29 b 3.98556915512e-06
R29 a 30 975.856685504
C29 30 b 3.39363842947e-06
R30 a 31 531.958176275
C30 31 b 2.8896203633e-06
R31 a 32 289.980593984
C31 32 b 2.46045830089e-06
R32 a 33 158.073977688
C32 33 b 2.09503474134e-06
R33 a 34 86.169153869
C33 34 b 1.78388333826e-06
R34 a 35 46.972456739
C34 35 b 1.51894367273e-06
R35 a 36 25.6055861411
C35 36 b 1.29335244713e-06
R36 a 37 13.9580955979
C36 37 b 1.10126569045e-06
R37 a 38 7.60882534167
C37 38 b 9.37707369436e-07
R38 a 39 4.14771647566
C38 39 b 7.98440483821e-07
R39 a 40 2.2609997194
C39 40 b 6.79857306217e-07
R40 a 41 1.23251426686
C40 41 b 5.78885923475e-07
R41 a 42 0.671867141321
C41 42 b 4.92910658358e-07
R42 a 43 0.366247651428
C42 43 b 4.19704310074e-07
R43 a 44 0.199648611946
C43 44 b 3.57370458332e-07
R44 a 45 0.108832283556
C44 45 b 3.0429433633e-07
R45 a 46 0.0593265629473
C45 46 b 2.59100999995e-07
R46 a 47 0.0323400461347
C46 47 b 2.20619709877e-07
R47 a 48 0.0176291787698
C47 48 b 1.87853602985e-07
R48 a 49 0.00961000311513
C48 49 b 1.59953868919e-07
R49 a 50 0.00523859682171
C49 50 b 1.36197761318e-07
R50 a 51 0.00285565949684
C50 51 b 1.15969875023e-07
R51 a 52 0.00155667470497
C51 52 b 9.8746203923e-08
R52 a 53 0.000848573206917
C52 53 b 8.40805665025e-08
R53 a 54 0.000462573513399
C53 54 b 7.15930474542e-08
R54 a 55 0.000252157684869
C54 55 b 6.09601559193e-08
R55 a b 10000000000.0
.ENDS displacement
****************************************
*          Combine subcircuits         *
****************************************
.SUBCKT interface a b
X_1 a n1 faradaic
X_2 a n1 displacement
R3 n1 b 13.38
.ENDS interface
****************************************
*          Circuit description         *
****************************************
X_ladder w1 w2 w3 w4 w5 w6 w7 w8 ladder
X_interface1 e1 w1 interface
X_interface2 e2 w2 interface
X_interface3 e3 w3 interface
X_interface4 e4 w4 interface
X_interface5 e5 w5 interface
X_interface6 e6 w6 interface
X_interface7 e7 w7 interface
X_interface8 e8 w8 interface
R_in 1 e7 0
R_out 0 e2 0
V1 1 0 DC 0 PWL(66 0.5 67 0.55 131 0.55 132 0.6 196 0.6 197 0.65 261 0.65 262 0.7 326 0.7 327 0.75 391 0.75 392 0.8 456 0.8 457 0.85 521 0.85 522 0.9 586 0.9 587 0.95 651 0.95 652 1.0 )
****************************************
*           Simulation options         *
****************************************
.control
TRAN 1 651 0
wrdata model_data v(e7,e2) i(V1) * -1.00 
.endc
.END
